/*
Let the two inputs be a[1:0] and b[1:0]. Then, the truth table would be 

| a[1] | a[0] | b[1] | b[0] | a_gt_b | 
|  0   |  0   |  0   |  0   |  0     | 
|  0   |  0   |  0   |  1   |  0     | 
|  0   |  0   |  1   |  0   |  0     | 
|  0   |  0   |  1   |  1   |  0     | 
|  0   |  1   |  0   |  0   |  1     | 
|  0   |  1   |  0   |  1   |  0     | 
|  0   |  1   |  1   |  0   |  0     | 
|  0   |  1   |  1   |  1   |  0     | 
|  1   |  0   |  0   |  0   |  1     | 
|  1   |  0   |  0   |  1   |  1     | 
|  1   |  0   |  1   |  0   |  0     | 
|  1   |  0   |  1   |  1   |  0     | 
|  1   |  1   |  0   |  0   |  1     | 
|  1   |  1   |  0   |  1   |  1     | 
|  1   |  1   |  1   |  0   |  1     | 
|  1   |  1   |  1   |  1   |  0     | 

a_gt_b = (a[1] . ~b[1]) + (a[1] . b[1] . a[0] . ~b[0]) + (~a[1] . ~b[1] . a[0] . ~b[0])
*/

module gt2 (
  input wire[1:0] a, b, 
  output wire a_gt_b
);

assign a_gt_b = (a[1] & ~b[1]) + (a[1] & b[1] & a[0] & ~b[0]) + (~a[1] & ~b[1] & a[0] & ~b[0]);
  
endmodule